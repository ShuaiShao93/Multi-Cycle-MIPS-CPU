module Bridge(
    input PClk,
    input IorD,
    input [31:2] PrA,
    input [3:0] PrBE,
    input [31:0] PrWData,
    output reg [31:0] PrRData,
    input PrReq,
    input PrRW,
    output reg PrReady,
    input [31:0] Din_IM,
    input [31:0] Din_DM,
    output reg [31:0] Dout_DM,
    output [12:2] A_IM,
    output [14:2] A_DM,
    output reg [3:0] BE,
    output reg We_DM,
    output [6:2] ADR_O, 
    output [7:0] DAT_O, 
    output reg WE_O, 
    input ACK_I_UART, 
    output STB_O_UART, 
    input [7:0] DAT_I_UART, 
    input ACK_I_TMR, 
    output reg STB_O_TMR, 
    input [7:0] DAT_I_TMR);
    `include "parameter.v"
    wire [1:0] aim;
    assign aim = (PrA[31:16] == 16'b1001000000000000)? AIM_DM :
               (PrA[31:14] == 18'b101111111100000000)? AIM_IM : AIM_WB;
    assign ADR_O = {PrA[10:8], PrA[3:2]};
    assign DAT_O = PrWData[7:0];
    assign A_IM = PrA[12:2];
    assign A_DM = PrA[14:2]; 
    always @(posedge PClk) begin
        if(PrReq)
            case(PrRW)
                RW_R:begin
                    if(aim == AIM_IM)
                      begin
                        PrRData[31:24] <= PrBE[3]? Din_IM[31:24] : 8'b0;
                        PrRData[23:16] <= PrBE[2]? Din_IM[23:16] : 8'b0;
                        PrRData[15:8]  <= PrBE[1]? Din_IM[15:8]  : 8'b0;
                        PrRData[7:0]   <= PrBE[0]? Din_IM[7:0]   : 8'b0;
                      end
                    else if(aim == AIM_DM)
                      begin
                        PrRData[31:24] <= PrBE[3]? Din_DM[31:24] : 8'b0;
                        PrRData[23:16] <= PrBE[2]? Din_DM[23:16] : 8'b0;
                        PrRData[15:8]  <= PrBE[1]? Din_DM[15:8]  : 8'b0;
                        PrRData[7:0]   <= PrBE[0]? Din_DM[7:0]   : 8'b0;
                      end
                    else if(aim == AIM_WB)
                      begin
                        PrRData[31:24] <= 8'b0;
                        PrRData[23:16] <= 8'b0;
                        PrRData[15:8] <= 8'b0;
                        PrRData[7:0] <= DAT_I_TMR;
                      end
                    PrReady <= 1;
                end
                RW_W: if(aim == AIM_DM)
                begin
                    Dout_DM[31:24] <= PrBE[3]? PrWData[31:24] : 8'b0;
                    Dout_DM[23:16] <= PrBE[2]? PrWData[23:16] : 8'b0;
                    Dout_DM[15:8]  <= PrBE[1]? PrWData[15:8] : 8'b0;
                    Dout_DM[7:0]   <= PrBE[0]? PrWData[7:0] : 8'b0;
                    PrReady <= 1;
                    BE <= PrBE;
                    We_DM <= 1;
                end
                else if(aim == AIM_WB)
                begin
                    WE_O <= 1;
                    STB_O_TMR <= 1;
                    PrReady <= 1;
                end
            endcase
        if(PrReady)
            PrReady <= 0;
        if(We_DM)
            We_DM <= 0;
        if(WE_O)
            WE_O <= 0;
    end
endmodule