module ALU(input [31:0] A, B, 
           input [4:0] Ctrl, 
           output reg [31:0] C, 
           output Zero, 
           output reg Compare);
    `include "parameter.v"
    always @(*)
        case (Ctrl)
            ALUOp_NOP : C <= B;
            ALUOp_ADDU : C <= A + B;
            ALUOp_ADD : C <= A + B;
            ALUOp_SUBU : C <= A - B;
            ALUOp_SUB : C <= A - B;
            ALUOp_AND : C <= A & B;
            ALUOp_OR : C <= A | B;
            ALUOp_NOR : C <= ~ (A | B);
            ALUOp_XOR : C <= A ^ B;
            ALUOp_SLTU : C <= (A < B)? 1 : 0;
            ALUOp_SLT : C <= ((A < B && A[31] == B[31]) || (A[31] > B[31]))? 1 : 0;
            ALUOp_LTZ : Compare <= (A[31] == 1)? 1 : 0;
            ALUOp_LEZ : Compare <= (A[31] == 1 ||  A == 0)? 1 : 0;
            ALUOp_GTZ : Compare <= (A[31] == 0 && A != 0)? 1 : 0;
            ALUOp_GEZ : Compare <= (A[31] == 0)? 1 : 0;
            ALUOp_SEQ : Compare <= (A == B)? 1 : 0;
            ALUOp_SNE : Compare <= (A != B)? 1 : 0;
    endcase
    assign Zero = (C == 0);
endmodule
